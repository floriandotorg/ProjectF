----------------------------------------------------------------------------------
-- company: 
-- engineer: 
-- 
-- create date:    18:42:25 05/21/2013 
-- design name: 
-- module name:    uart - behavioral 
-- project name: 
-- target devices: 
-- tool versions: 
-- description: 
--
-- dependencies: 
--
-- revision: 
-- revision 0.01 - file created
-- additional comments: 
--
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

-- uncomment the following library declaration if using
-- arithmetic functions with signed or unsigned values
--use ieee.numeric_std.all;

-- uncomment the following library declaration if instantiating
-- any xilinx primitives in this code.
--library unisim;
--use unisim.vcomponents.all;

entity uart is
    port ( clk : in  std_logic );
end uart;

architecture behavioral of uart is

begin


end behavioral;

